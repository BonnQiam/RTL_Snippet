//----------------------------------------------------
//（参数化）n-m 译码器
// a：输入为二进制数（宽度为 n）
// b：输出为独热码（宽度为 m）
//-----------------------------------------------------
module Dec_n_m (
    a,b
);
    parameter n = 2;//设置默认值
    parameter m = 4;

    input   [n-1:0] a;
    output  [m-1:0] b;

    assign b = 1 << a; 
    /*
        采用左移运算符 "<<" ，根据输入 a 将 1 移动到指定位置，
        并且以独热码的形式将结果从 b 输出
    */
endmodule
